Voltage divider circuit

V1 Vin 0 5V
R1 Vin Vout 1k
R2 Vout 0 2k

* Does not work with Ngspice
* .step param R 1k 5k 1k

.tran 100m 1
.op
.end 


