**.subckt inv_tran
Vin Vin GND pulse(0 1.8 0 1ns 1ns 4ns 10ns)
Vdd Vdd GND 1.8
x1 Vdd Vout Vin GND inv_1
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt



.include /home/harshit/.xschem/inv.spice
.tran 100ps 20ns
.save all
.end

**** end user architecture code
**.ends

* expanding   symbol:  /home/harshit/.xschem/inv_1.sym # of pins=4
* sym_path: /home/harshit/.xschem/inv_1.sym
* sch_path: /home/harshit/.xschem/inv_1.sch
.subckt inv_1  Vdd Vout Vin VSS
*.ipin Vdd
*.ipin VSS
*.opin Vout
*.ipin Vin
XM1 Vout Vin VSS VSS sky130_fd_pr__nfet_01v8 L=0.30 W=3.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vout Vin Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.30 W=3.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
